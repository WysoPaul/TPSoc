// SysHdwTP.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module SysHdwTP (
		input  wire        bp1_export,    //   bp1.export
		input  wire        clk_clk,       //   clk.clk
		input  wire        reset_reset_n, // reset.reset_n
		output wire [47:0] s7seg_export   // s7seg.export
	);

	wire  [31:0] nios_data_master_readdata;                            // mm_interconnect_0:NIOS_data_master_readdata -> NIOS:d_readdata
	wire         nios_data_master_waitrequest;                         // mm_interconnect_0:NIOS_data_master_waitrequest -> NIOS:d_waitrequest
	wire         nios_data_master_debugaccess;                         // NIOS:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NIOS_data_master_debugaccess
	wire  [17:0] nios_data_master_address;                             // NIOS:d_address -> mm_interconnect_0:NIOS_data_master_address
	wire   [3:0] nios_data_master_byteenable;                          // NIOS:d_byteenable -> mm_interconnect_0:NIOS_data_master_byteenable
	wire         nios_data_master_read;                                // NIOS:d_read -> mm_interconnect_0:NIOS_data_master_read
	wire         nios_data_master_readdatavalid;                       // mm_interconnect_0:NIOS_data_master_readdatavalid -> NIOS:d_readdatavalid
	wire         nios_data_master_write;                               // NIOS:d_write -> mm_interconnect_0:NIOS_data_master_write
	wire  [31:0] nios_data_master_writedata;                           // NIOS:d_writedata -> mm_interconnect_0:NIOS_data_master_writedata
	wire  [31:0] nios_instruction_master_readdata;                     // mm_interconnect_0:NIOS_instruction_master_readdata -> NIOS:i_readdata
	wire         nios_instruction_master_waitrequest;                  // mm_interconnect_0:NIOS_instruction_master_waitrequest -> NIOS:i_waitrequest
	wire  [17:0] nios_instruction_master_address;                      // NIOS:i_address -> mm_interconnect_0:NIOS_instruction_master_address
	wire         nios_instruction_master_read;                         // NIOS:i_read -> mm_interconnect_0:NIOS_instruction_master_read
	wire         nios_instruction_master_readdatavalid;                // mm_interconnect_0:NIOS_instruction_master_readdatavalid -> NIOS:i_readdatavalid
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;  // mm_interconnect_0:JTAG_avalon_jtag_slave_chipselect -> JTAG:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;    // JTAG:av_readdata -> mm_interconnect_0:JTAG_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest; // JTAG:av_waitrequest -> mm_interconnect_0:JTAG_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;     // mm_interconnect_0:JTAG_avalon_jtag_slave_address -> JTAG:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;        // mm_interconnect_0:JTAG_avalon_jtag_slave_read -> JTAG:av_read_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;       // mm_interconnect_0:JTAG_avalon_jtag_slave_write -> JTAG:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;   // mm_interconnect_0:JTAG_avalon_jtag_slave_writedata -> JTAG:av_writedata
	wire  [31:0] mm_interconnect_0_nios_debug_mem_slave_readdata;      // NIOS:debug_mem_slave_readdata -> mm_interconnect_0:NIOS_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios_debug_mem_slave_waitrequest;   // NIOS:debug_mem_slave_waitrequest -> mm_interconnect_0:NIOS_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios_debug_mem_slave_debugaccess;   // mm_interconnect_0:NIOS_debug_mem_slave_debugaccess -> NIOS:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios_debug_mem_slave_address;       // mm_interconnect_0:NIOS_debug_mem_slave_address -> NIOS:debug_mem_slave_address
	wire         mm_interconnect_0_nios_debug_mem_slave_read;          // mm_interconnect_0:NIOS_debug_mem_slave_read -> NIOS:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios_debug_mem_slave_byteenable;    // mm_interconnect_0:NIOS_debug_mem_slave_byteenable -> NIOS:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios_debug_mem_slave_write;         // mm_interconnect_0:NIOS_debug_mem_slave_write -> NIOS:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios_debug_mem_slave_writedata;     // mm_interconnect_0:NIOS_debug_mem_slave_writedata -> NIOS:debug_mem_slave_writedata
	wire         mm_interconnect_0_memoire_s1_chipselect;              // mm_interconnect_0:MEMOIRE_s1_chipselect -> MEMOIRE:chipselect
	wire  [31:0] mm_interconnect_0_memoire_s1_readdata;                // MEMOIRE:readdata -> mm_interconnect_0:MEMOIRE_s1_readdata
	wire  [13:0] mm_interconnect_0_memoire_s1_address;                 // mm_interconnect_0:MEMOIRE_s1_address -> MEMOIRE:address
	wire   [3:0] mm_interconnect_0_memoire_s1_byteenable;              // mm_interconnect_0:MEMOIRE_s1_byteenable -> MEMOIRE:byteenable
	wire         mm_interconnect_0_memoire_s1_write;                   // mm_interconnect_0:MEMOIRE_s1_write -> MEMOIRE:write
	wire  [31:0] mm_interconnect_0_memoire_s1_writedata;               // mm_interconnect_0:MEMOIRE_s1_writedata -> MEMOIRE:writedata
	wire         mm_interconnect_0_memoire_s1_clken;                   // mm_interconnect_0:MEMOIRE_s1_clken -> MEMOIRE:clken
	wire   [7:0] mm_interconnect_0_ip7seg_s1_readdata;                 // IP7Seg:avs_s1_readdata -> mm_interconnect_0:IP7Seg_s1_readdata
	wire   [2:0] mm_interconnect_0_ip7seg_s1_address;                  // mm_interconnect_0:IP7Seg_s1_address -> IP7Seg:avs_s1_address
	wire         mm_interconnect_0_ip7seg_s1_read;                     // mm_interconnect_0:IP7Seg_s1_read -> IP7Seg:avs_s1_read
	wire         mm_interconnect_0_ip7seg_s1_write;                    // mm_interconnect_0:IP7Seg_s1_write -> IP7Seg:avs_s1_write
	wire   [7:0] mm_interconnect_0_ip7seg_s1_writedata;                // mm_interconnect_0:IP7Seg_s1_writedata -> IP7Seg:avs_s1_writedata
	wire         mm_interconnect_0_ip_bp1_s1_chipselect;               // mm_interconnect_0:IP_BP1_s1_chipselect -> IP_BP1:chipselect
	wire  [31:0] mm_interconnect_0_ip_bp1_s1_readdata;                 // IP_BP1:readdata -> mm_interconnect_0:IP_BP1_s1_readdata
	wire   [1:0] mm_interconnect_0_ip_bp1_s1_address;                  // mm_interconnect_0:IP_BP1_s1_address -> IP_BP1:address
	wire         mm_interconnect_0_ip_bp1_s1_write;                    // mm_interconnect_0:IP_BP1_s1_write -> IP_BP1:write_n
	wire  [31:0] mm_interconnect_0_ip_bp1_s1_writedata;                // mm_interconnect_0:IP_BP1_s1_writedata -> IP_BP1:writedata
	wire         irq_mapper_receiver0_irq;                             // JTAG:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                             // IP_BP1:irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios_irq_irq;                                         // irq_mapper:sender_irq -> NIOS:irq
	wire         rst_controller_reset_out_reset;                       // rst_controller:reset_out -> [IP7Seg:avs_s1_reset, IP_BP1:reset_n, JTAG:rst_n, MEMOIRE:reset, NIOS:reset_n, irq_mapper:reset, mm_interconnect_0:NIOS_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                   // rst_controller:reset_req -> [MEMOIRE:reset_req, NIOS:reset_req, rst_translator:reset_req_in]
	wire         nios_debug_reset_request_reset;                       // NIOS:debug_reset_request -> rst_controller:reset_in1

	seg7_if #(
		.SEG7_NUM       (6),
		.ADDR_WIDTH     (3),
		.DEFAULT_ACTIVE (1),
		.LOW_ACTIVE     (1)
	) ip7seg (
		.avs_s1_clk         (clk_clk),                               //       s1_clock.clk
		.avs_s1_reset       (rst_controller_reset_out_reset),        // s1_clock_reset.reset
		.avs_s1_address     (mm_interconnect_0_ip7seg_s1_address),   //             s1.address
		.avs_s1_read        (mm_interconnect_0_ip7seg_s1_read),      //               .read
		.avs_s1_readdata    (mm_interconnect_0_ip7seg_s1_readdata),  //               .readdata
		.avs_s1_write       (mm_interconnect_0_ip7seg_s1_write),     //               .write
		.avs_s1_writedata   (mm_interconnect_0_ip7seg_s1_writedata), //               .writedata
		.avs_s1_export_seg7 (s7seg_export)                           //      s1_export.export
	);

	SysHdwTP_IP_BP1 ip_bp1 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_ip_bp1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ip_bp1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ip_bp1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ip_bp1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ip_bp1_s1_readdata),   //                    .readdata
		.in_port    (bp1_export),                             // external_connection.export
		.irq        (irq_mapper_receiver1_irq)                //                 irq.irq
	);

	SysHdwTP_JTAG jtag (
		.clk            (clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                              //               irq.irq
	);

	SysHdwTP_MEMOIRE memoire (
		.clk        (clk_clk),                                 //   clk1.clk
		.address    (mm_interconnect_0_memoire_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_memoire_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_memoire_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_memoire_s1_write),      //       .write
		.readdata   (mm_interconnect_0_memoire_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_memoire_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_memoire_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),          // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),      //       .reset_req
		.freeze     (1'b0)                                     // (terminated)
	);

	SysHdwTP_NIOS nios (
		.clk                                 (clk_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                    //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                 //                          .reset_req
		.d_address                           (nios_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios_data_master_read),                              //                          .read
		.d_readdata                          (nios_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios_data_master_write),                             //                          .write
		.d_writedata                         (nios_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios_instruction_master_read),                       //                          .read
		.i_readdata                          (nios_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                    // custom_instruction_master.readra
	);

	SysHdwTP_mm_interconnect_0 mm_interconnect_0 (
		.CLOCK_clk_clk                          (clk_clk),                                              //                        CLOCK_clk.clk
		.NIOS_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                       // NIOS_reset_reset_bridge_in_reset.reset
		.NIOS_data_master_address               (nios_data_master_address),                             //                 NIOS_data_master.address
		.NIOS_data_master_waitrequest           (nios_data_master_waitrequest),                         //                                 .waitrequest
		.NIOS_data_master_byteenable            (nios_data_master_byteenable),                          //                                 .byteenable
		.NIOS_data_master_read                  (nios_data_master_read),                                //                                 .read
		.NIOS_data_master_readdata              (nios_data_master_readdata),                            //                                 .readdata
		.NIOS_data_master_readdatavalid         (nios_data_master_readdatavalid),                       //                                 .readdatavalid
		.NIOS_data_master_write                 (nios_data_master_write),                               //                                 .write
		.NIOS_data_master_writedata             (nios_data_master_writedata),                           //                                 .writedata
		.NIOS_data_master_debugaccess           (nios_data_master_debugaccess),                         //                                 .debugaccess
		.NIOS_instruction_master_address        (nios_instruction_master_address),                      //          NIOS_instruction_master.address
		.NIOS_instruction_master_waitrequest    (nios_instruction_master_waitrequest),                  //                                 .waitrequest
		.NIOS_instruction_master_read           (nios_instruction_master_read),                         //                                 .read
		.NIOS_instruction_master_readdata       (nios_instruction_master_readdata),                     //                                 .readdata
		.NIOS_instruction_master_readdatavalid  (nios_instruction_master_readdatavalid),                //                                 .readdatavalid
		.IP7Seg_s1_address                      (mm_interconnect_0_ip7seg_s1_address),                  //                        IP7Seg_s1.address
		.IP7Seg_s1_write                        (mm_interconnect_0_ip7seg_s1_write),                    //                                 .write
		.IP7Seg_s1_read                         (mm_interconnect_0_ip7seg_s1_read),                     //                                 .read
		.IP7Seg_s1_readdata                     (mm_interconnect_0_ip7seg_s1_readdata),                 //                                 .readdata
		.IP7Seg_s1_writedata                    (mm_interconnect_0_ip7seg_s1_writedata),                //                                 .writedata
		.IP_BP1_s1_address                      (mm_interconnect_0_ip_bp1_s1_address),                  //                        IP_BP1_s1.address
		.IP_BP1_s1_write                        (mm_interconnect_0_ip_bp1_s1_write),                    //                                 .write
		.IP_BP1_s1_readdata                     (mm_interconnect_0_ip_bp1_s1_readdata),                 //                                 .readdata
		.IP_BP1_s1_writedata                    (mm_interconnect_0_ip_bp1_s1_writedata),                //                                 .writedata
		.IP_BP1_s1_chipselect                   (mm_interconnect_0_ip_bp1_s1_chipselect),               //                                 .chipselect
		.JTAG_avalon_jtag_slave_address         (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //           JTAG_avalon_jtag_slave.address
		.JTAG_avalon_jtag_slave_write           (mm_interconnect_0_jtag_avalon_jtag_slave_write),       //                                 .write
		.JTAG_avalon_jtag_slave_read            (mm_interconnect_0_jtag_avalon_jtag_slave_read),        //                                 .read
		.JTAG_avalon_jtag_slave_readdata        (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                                 .readdata
		.JTAG_avalon_jtag_slave_writedata       (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                                 .writedata
		.JTAG_avalon_jtag_slave_waitrequest     (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                                 .waitrequest
		.JTAG_avalon_jtag_slave_chipselect      (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  //                                 .chipselect
		.MEMOIRE_s1_address                     (mm_interconnect_0_memoire_s1_address),                 //                       MEMOIRE_s1.address
		.MEMOIRE_s1_write                       (mm_interconnect_0_memoire_s1_write),                   //                                 .write
		.MEMOIRE_s1_readdata                    (mm_interconnect_0_memoire_s1_readdata),                //                                 .readdata
		.MEMOIRE_s1_writedata                   (mm_interconnect_0_memoire_s1_writedata),               //                                 .writedata
		.MEMOIRE_s1_byteenable                  (mm_interconnect_0_memoire_s1_byteenable),              //                                 .byteenable
		.MEMOIRE_s1_chipselect                  (mm_interconnect_0_memoire_s1_chipselect),              //                                 .chipselect
		.MEMOIRE_s1_clken                       (mm_interconnect_0_memoire_s1_clken),                   //                                 .clken
		.NIOS_debug_mem_slave_address           (mm_interconnect_0_nios_debug_mem_slave_address),       //             NIOS_debug_mem_slave.address
		.NIOS_debug_mem_slave_write             (mm_interconnect_0_nios_debug_mem_slave_write),         //                                 .write
		.NIOS_debug_mem_slave_read              (mm_interconnect_0_nios_debug_mem_slave_read),          //                                 .read
		.NIOS_debug_mem_slave_readdata          (mm_interconnect_0_nios_debug_mem_slave_readdata),      //                                 .readdata
		.NIOS_debug_mem_slave_writedata         (mm_interconnect_0_nios_debug_mem_slave_writedata),     //                                 .writedata
		.NIOS_debug_mem_slave_byteenable        (mm_interconnect_0_nios_debug_mem_slave_byteenable),    //                                 .byteenable
		.NIOS_debug_mem_slave_waitrequest       (mm_interconnect_0_nios_debug_mem_slave_waitrequest),   //                                 .waitrequest
		.NIOS_debug_mem_slave_debugaccess       (mm_interconnect_0_nios_debug_mem_slave_debugaccess)    //                                 .debugaccess
	);

	SysHdwTP_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios_irq_irq)                    //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios_debug_reset_request_reset),     // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
