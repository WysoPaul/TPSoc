
module SysHdwTP (
	bp1_export,
	clk_clk,
	reset_reset_n,
	s7seg_export);	

	input		bp1_export;
	input		clk_clk;
	input		reset_reset_n;
	output	[47:0]	s7seg_export;
endmodule
